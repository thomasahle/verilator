// Package that includes the class file
package DriverPkg;
   `include "DriverProxy.sv"
endpackage
