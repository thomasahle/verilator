// Minimal UVM package stub for testing assertions
package uvm_pkg;
  typedef enum {UVM_NONE=0, UVM_LOW=100, UVM_MEDIUM=200, UVM_HIGH=300, UVM_FULL=400, UVM_DEBUG=500} uvm_verbosity;
endpackage
