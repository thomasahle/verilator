// DESCRIPTION: Verilator: Test I2S AVIP
// Wrapper module that instantiates hdlTop and hvlTop from I2S AVIP
module tb_top;
  hdlTop hdl();
  hvlTop hvl();
endmodule
